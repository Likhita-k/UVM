class adder_sqr extends uvm_sequencer#(adder_tx);
`uvm_component_utils(adder_sqr)
`NEW_COMPONENT
endclass
