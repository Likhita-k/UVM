`define NUM 8

`include "uvm_pkg.sv"
import uvm_pkg::*;

`include "adder.v"
`include "common.sv"
`include "tx.sv"
`include "seq.sv"
`include "scb.sv"
`include "mon.sv"
`include "drv.sv"
`include "sqr.sv"
`include "agent.sv"
`include "env.sv"
`include "intf.sv"
`include "test_lib.sv"
`include "top.sv"
